module ejercicio_21(
    
    input A, B, C,
    output Y
);
    assign Y = !A;
endmodule